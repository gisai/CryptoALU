----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/18/2021 07:24:48 PM
-- Design Name: 
-- Module Name: extSigno - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Extensor_De_Signo is
    Port ( inmed : in STD_LOGIC_VECTOR (15 downto 0);
           salida : inout STD_LOGIC_VECTOR (31 downto 0));
end Extensor_De_Signo;

architecture Behavioral of Extensor_De_Signo is

begin

salida <= x"0000" & inmed when inmed(15)='0' ELSE
          x"FFFF" & inmed when inmed(15)='1';

end Behavioral;
